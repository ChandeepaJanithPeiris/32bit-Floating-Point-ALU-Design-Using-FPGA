library verilog;
use verilog.vl_types.all;
entity binary_div_tb is
end binary_div_tb;
