library verilog;
use verilog.vl_types.all;
entity binary_multiplier_tb is
end binary_multiplier_tb;
