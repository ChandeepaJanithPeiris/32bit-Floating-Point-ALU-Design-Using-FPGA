library verilog;
use verilog.vl_types.all;
entity fp_multiplier_tb is
end fp_multiplier_tb;
