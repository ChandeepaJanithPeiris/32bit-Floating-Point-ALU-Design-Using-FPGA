module binary_division (
    input logic [23:0] Q, // 24-bit dividend
    input logic [23:0] M, // 24-bit divisor
    output logic signed [24:0] Qo,  // 25-bit quotient
    output logic signed [24:0] A   // 25-bit remainder
);

logic signed [24:0] M_extended;
logic signed [24:0] A_new;
logic [23:0] Q_local;



always_comb begin
    A = 25'b0;  // Initialize A to zero
    M_extended = {1'b0, M};  // Extend M to 25 bits
    Q_local = Q;  // Local copy of Q
    Qo = 25'b0;  // Initialize Qo

    for (int i = 24; i > 0; i--) begin
        // Shift left A and Q
        A = {A[23:0], Q_local[23]};  
        Q_local = Q_local << 1;

        // Subtract M_extended from A
        A_new = A - M_extended;

        // Check if subtraction result is negative
        if (A_new[24] == 1) begin
            Qo = {Qo[23:0], 1'b0};  // Append 0 to Qo
        end
        else begin
            Qo = {Qo[23:0], 1'b1};  // Append 1 to Qo
            A = A_new;  // Update A with the new value
        end
    end
end

endmodule
