library verilog;
use verilog.vl_types.all;
entity extended_div_tb is
end extended_div_tb;
