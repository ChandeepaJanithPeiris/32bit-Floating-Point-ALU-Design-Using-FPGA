library verilog;
use verilog.vl_types.all;
entity binary_division_tb is
end binary_division_tb;
