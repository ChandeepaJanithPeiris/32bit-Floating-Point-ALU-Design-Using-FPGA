library verilog;
use verilog.vl_types.all;
entity right_shift_tb is
end right_shift_tb;
