module binary_multiplier #(parameter N = 24) (
    input  logic [N-1:0] A,  // N-bit input A
    input  logic [N-1:0] B,  // N-bit input B
    output logic [2*N-1:0] P // 2N-bit product
);

    // Array to hold partial products
    logic [2*N-1:0] partial_products [N-1:0];
    
    // Generate Partial Products using a generate block with genvar
    genvar i;
    generate
        for (i = 0; i < N; i = i + 1) begin : gen_partial_products
            assign partial_products[i] = (A & {N{B[i]}}) << i;
        end
    endgenerate

    // Sum up the partial products using an always block
    always_comb begin
        P = partial_products[0];  // Initialize sum with the first partial product
        for (int j = 1; j < N; j = j + 1) begin
            P = P + partial_products[j];  // Sum the partial products
        end
    end

endmodule
