library verilog;
use verilog.vl_types.all;
entity fp_adder_tb is
end fp_adder_tb;
