library verilog;
use verilog.vl_types.all;
entity fp_division_tb is
end fp_division_tb;
